package pack_util is
	constant NBREG: natural := 8
	type 

  
end package pack_util;

-- Package Body Section
package body pack_util is

end package body pack_util;